`ifndef ACX_BUILD_TIMESTAMP
`define ACX_BUILD_TIMESTAMP 32'h10201021
`endif
