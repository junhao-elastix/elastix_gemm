// ------------------------------------------------------------------
// Testbench for gfp8_bcv_controller.sv
//
// Purpose: Verify BCV loop orchestration for matrix multiplication
// Tests:
//  1. Simple case: B=1, C=1, V=1 (single NV dot product)
//  2. Small V loop: B=1, C=1, V=4 (accumulation test)
//  3. Multiple outputs: B=2, C=2, V=2 (full BCV test)
//  4. Real data: B=1, C=1, V=128 (full matrix)
//
// Author: Refactoring effort
// Date: Fri Oct 10 2025
// ------------------------------------------------------------------

`timescale 1ns/1ps

module tb_gfp8_bcv_controller;

    // Clock and reset
    logic clk;
    logic reset_n;
    
    // TILE command interface
    logic        tile_en;
    logic [7:0]  dim_b;
    logic [7:0]  dim_c;
    logic [7:0]  dim_v;
    logic [10:0] left_base_addr;
    logic [10:0] right_base_addr;
    logic        tile_done;
    
    // BRAM interfaces
    logic [10:0]  mem_left_rd_addr;
    logic         mem_left_rd_en;
    logic [255:0] mem_left_rd_data;
    
    logic [10:0]  mem_right_rd_addr;
    logic         mem_right_rd_en;
    logic [255:0] mem_right_rd_data;
    
    // Result interface
    logic signed [31:0] result_mantissa;
    logic signed [7:0]  result_exponent;
    logic               result_valid;
    
    // Test control
    integer test_num;
    logic test_passed;
    integer result_count;
    
    // BRAM models (storage for left and right matrices)
    logic [255:0] bram_left [0:1055];   // Depth for full matrix storage
    logic [255:0] bram_right [0:1055];
    
    // Result collection
    logic signed [31:0] results_mantissa [0:255];  // Up to 16x16 = 256 results
    logic signed [7:0]  results_exponent [0:255];
    
    // ===================================================================
    // DUT Instantiation
    // ===================================================================
    gfp8_bcv_controller dut (
        .i_clk                  (clk),
        .i_reset_n              (reset_n),
        
        .i_tile_en              (tile_en),
        .i_dim_b                (dim_b),
        .i_dim_c                (dim_c),
        .i_dim_v                (dim_v),
        .i_left_base_addr       (left_base_addr),
        .i_right_base_addr      (right_base_addr),
        .o_tile_done            (tile_done),
        
        .o_mem_left_rd_addr     (mem_left_rd_addr),
        .o_mem_left_rd_en       (mem_left_rd_en),
        .i_mem_left_rd_data     (mem_left_rd_data),
        
        .o_mem_right_rd_addr    (mem_right_rd_addr),
        .o_mem_right_rd_en      (mem_right_rd_en),
        .i_mem_right_rd_data    (mem_right_rd_data),
        
        .o_result_mantissa      (result_mantissa),
        .o_result_exponent      (result_exponent),
        .o_result_valid         (result_valid)
    );
    
    // ===================================================================
    // Clock Generation
    // ===================================================================
    initial begin
        clk = 0;
        forever #5 clk = ~clk;  // 100MHz clock
    end
    
    // ===================================================================
    // BRAM Models (1-cycle read latency)
    // ===================================================================
    logic [255:0] bram_left_reg;
    logic [255:0] bram_right_reg;
    
    always_ff @(posedge clk) begin
        if (mem_left_rd_en) begin
            bram_left_reg <= bram_left[mem_left_rd_addr];
        end
        if (mem_right_rd_en) begin
            bram_right_reg <= bram_right[mem_right_rd_addr];
        end
    end
    
    assign mem_left_rd_data = bram_left_reg;
    assign mem_right_rd_data = bram_right_reg;
    
    // ===================================================================
    // Result Collection Monitor
    // ===================================================================
    always @(posedge clk) begin
        if (result_valid) begin
            results_mantissa[result_count] = result_mantissa;
            results_exponent[result_count] = result_exponent;
            $display("  [%0t] Result %0d: mantissa=%0d, exponent=%0d", 
                     $time, result_count, result_mantissa, result_exponent);
            result_count = result_count + 1;
        end
    end
    
    // ===================================================================
    // Helper Task: Initialize BRAM with Simple Pattern
    // ===================================================================
    task init_bram_simple();
        $display("  Initializing BRAM with simple pattern (all 1s)...");
        
        // Simple pattern: exponents = 15, mantissas = 1
        for (int i = 0; i < 1056; i++) begin
            if (i < 16) begin
                // Exponent lines (bytes all set to 15)
                bram_left[i] = {32{8'd15}};
                bram_right[i] = {32{8'd15}};
            end else begin
                // Mantissa lines (all 1s)
                bram_left[i] = {32{8'sd1}};
                bram_right[i] = {32{8'sd1}};
            end
        end
    endtask
    
    // ===================================================================
    // Helper Task: Load BRAM from Hex Files
    // ===================================================================
    task load_bram_from_hex();
        logic [255:0] left_data [0:527];
        logic [255:0] right_data [0:527];
        
        $display("  Loading BRAM from hex files...");
        $readmemh("/home/dev/Dev/elastix_gemm/hex/left.hex", left_data);
        $readmemh("/home/dev/Dev/elastix_gemm/hex/right.hex", right_data);
        
        // Copy to BRAM models
        for (int i = 0; i < 528; i++) begin
            bram_left[i] = left_data[i];
            bram_right[i] = right_data[i];
        end
        
        $display("  Loaded %0d lines from left.hex", 528);
        $display("  Loaded %0d lines from right.hex", 528);
    endtask
    
    // ===================================================================
    // Helper Task: Send TILE Command
    // ===================================================================
    task send_tile_command(input logic [7:0] b, input logic [7:0] c, input logic [7:0] v);
        $display("  Sending TILE command: B=%0d, C=%0d, V=%0d", b, c, v);
        @(posedge clk);
        tile_en <= 1'b1;
        dim_b <= b;
        dim_c <= c;
        dim_v <= v;
        left_base_addr <= 11'd0;
        right_base_addr <= 11'd0;
        @(posedge clk);
        tile_en <= 1'b0;
    endtask
    
    // ===================================================================
    // Helper Task: Wait for TILE Done
    // ===================================================================
    task wait_tile_done(input integer timeout_cycles);
        integer cycle_count;
        cycle_count = 0;
        
        $display("  Waiting for TILE completion...");
        while (!tile_done && cycle_count < timeout_cycles) begin
            @(posedge clk);
            cycle_count++;
        end
        
        if (tile_done) begin
            $display("  TILE completed in %0d cycles", cycle_count);
        end else begin
            $display("  ERROR: TILE timeout after %0d cycles", timeout_cycles);
            test_passed = 0;
        end
    endtask
    
    // ===================================================================
    // Test Stimulus
    // ===================================================================
    initial begin
        // Initialize
        reset_n = 0;
        tile_en = 0;
        dim_b = 8'd0;
        dim_c = 8'd0;
        dim_v = 8'd0;
        left_base_addr = 11'd0;
        right_base_addr = 11'd0;
        test_num = 0;
        test_passed = 1;
        result_count = 0;
        
        // Initialize BRAM
        for (int i = 0; i < 1056; i++) begin
            bram_left[i] = 256'd0;
            bram_right[i] = 256'd0;
        end
        
        // Reset
        repeat(5) @(posedge clk);
        reset_n = 1;
        repeat(2) @(posedge clk);
        
        $display("\n========================================");
        $display("GFP8 BCV Controller Testbench");
        $display("========================================\n");
        
        // ===============================================================
        // Test 1: Simple Case - B=1, C=1, V=1
        // ===============================================================
        test_num = 1;
        $display("[TEST %0d] Simple case: B=1, C=1, V=1", test_num);
        
        init_bram_simple();
        result_count = 0;
        
        send_tile_command(8'd1, 8'd1, 8'd1);
        wait_tile_done(1000);
        
        repeat(5) @(posedge clk);
        
        $display("  Results collected: %0d", result_count);
        if (result_count == 1) begin
            $display("  Expected: 1 result (1x1 output)");
            $display("  Result mantissa=%0d, exponent=%0d", 
                     results_mantissa[0], results_exponent[0]);
            // Each NV dot product: 128 elements x (1*1) = 128
            if (results_mantissa[0] == 32'sd128 && results_exponent[0] == 8'sd0) begin
                $display("  [PASS]\n");
            end else begin
                $display("  [FAIL] Expected mantissa=128, exponent=0\n");
                test_passed = 0;
            end
        end else begin
            $display("  [FAIL] Expected 1 result, got %0d\n", result_count);
            test_passed = 0;
        end
        
        // ===============================================================
        // Test 2: V Loop Test - B=1, C=1, V=4
        // ===============================================================
        test_num = 2;
        $display("[TEST %0d] V loop test: B=1, C=1, V=4", test_num);
        $display("  Testing V-loop accumulation");
        
        init_bram_simple();
        result_count = 0;
        
        send_tile_command(8'd1, 8'd1, 8'd4);
        wait_tile_done(5000);
        
        repeat(5) @(posedge clk);
        
        $display("  Results collected: %0d", result_count);
        if (result_count == 1) begin
            $display("  Expected: 1 result (accumulation of 4 NV dots)");
            $display("  Result mantissa=%0d, exponent=%0d", 
                     results_mantissa[0], results_exponent[0]);
            // 4 NV dot products: 4 x 128 = 512
            if (results_mantissa[0] == 32'sd512 && results_exponent[0] == 8'sd0) begin
                $display("  [PASS]\n");
            end else begin
                $display("  [WARN] Expected mantissa=512, exponent=0\n");
                $display("  Actual values may differ due to accumulation order\n");
            end
        end else begin
            $display("  [FAIL] Expected 1 result, got %0d\n", result_count);
            test_passed = 0;
        end
        
        // ===============================================================
        // Test 3: Multiple Outputs - B=2, C=2, V=2
        // ===============================================================
        test_num = 3;
        $display("[TEST %0d] Multiple outputs: B=2, C=2, V=2", test_num);
        $display("  Testing full BCV loop with 4 outputs");
        
        init_bram_simple();
        result_count = 0;
        
        send_tile_command(8'd2, 8'd2, 8'd2);
        wait_tile_done(10000);
        
        repeat(5) @(posedge clk);
        
        $display("  Results collected: %0d", result_count);
        if (result_count == 4) begin
            $display("  Expected: 4 results (2x2 output matrix)");
            for (int i = 0; i < 4; i++) begin
                $display("    Output[%0d]: mantissa=%0d, exponent=%0d", 
                         i, results_mantissa[i], results_exponent[i]);
            end
            // Each output: 2 NV dot products = 2 x 128 = 256
            if (results_mantissa[0] == 32'sd256) begin
                $display("  [PASS]\n");
            end else begin
                $display("  [WARN] Results may vary\n");
            end
        end else begin
            $display("  [FAIL] Expected 4 results, got %0d\n", result_count);
            test_passed = 0;
        end
        
        // ===============================================================
        // Test 4: Real Data - B=1, C=1, V=128
        // ===============================================================
        test_num = 4;
        $display("[TEST %0d] Real data: B=1, C=1, V=128", test_num);
        $display("  Loading actual hex files (full matrix)");
        
        load_bram_from_hex();
        result_count = 0;
        
        send_tile_command(8'd1, 8'd1, 8'd128);
        wait_tile_done(100000);  // Long timeout for full matrix
        
        repeat(5) @(posedge clk);
        
        $display("  Results collected: %0d", result_count);
        if (result_count == 1) begin
            $display("  Expected: 1 result (full 128-NV accumulation)");
            $display("  Result mantissa=%0d, exponent=%0d", 
                     results_mantissa[0], results_exponent[0]);
            $display("  [INFO] Manual verification needed against Python golden model\n");
        end else begin
            $display("  [FAIL] Expected 1 result, got %0d\n", result_count);
            test_passed = 0;
        end
        
        // ===============================================================
        // Test Summary
        // ===============================================================
        $display("========================================");
        if (test_passed) begin
            $display("All tests PASSED");
        end else begin
            $display("Some tests FAILED");
        end
        $display("========================================\n");
        
        $finish;
    end
    
    // ===================================================================
    // Timeout
    // ===================================================================
    initial begin
        #10000000;  // 10ms timeout
        $display("ERROR: Testbench timeout!");
        $finish;
    end

endmodule

