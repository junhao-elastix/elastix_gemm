// ------------------------------------------------------------------
// Testbench for GFP8 Group Dot Product Module
//
// Purpose: Validate 32-pair GFP8 dot product computation
// Test Cases:
//  1. First group from left.hex and right.hex
//  2. Zero exponent handling
//  3. Known values with manual calculation
//
// Author: Refactoring verification
// Date: Thu Oct 9 2025
// ------------------------------------------------------------------

`timescale 1ns/1ps

module tb_gfp8_group_dot;

    // ===================================================================
    // Testbench Signals
    // ===================================================================
    logic         clk;
    logic         reset_n;
    
    logic [4:0]   exp_left;
    logic [255:0] man_left;
    logic [4:0]   exp_right;
    logic [255:0] man_right;
    
    logic signed [31:0] result_mantissa;
    logic signed [7:0]  result_exponent;
    
    // ===================================================================
    // Clock Generation (100 MHz)
    // ===================================================================
    initial begin
        clk = 0;
        forever #5 clk = ~clk;  // 10ns period = 100MHz
    end
    
    // ===================================================================
    // DUT Instantiation
    // ===================================================================
    gfp8_group_dot_mlp dut (
        .i_clk              (clk),
        .i_reset_n          (reset_n),
        .i_exp_left         (exp_left),
        .i_man_left         (man_left),
        .i_exp_right        (exp_right),
        .i_man_right        (man_right),
        .o_result_mantissa  (result_mantissa),
        .o_result_exponent  (result_exponent)
    );
    
    // ===================================================================
    // Helper Functions
    // ===================================================================
    
    // Display result in readable format
    task display_result(input string test_name);
        real fp_value;
        
        // Calculate floating-point value: mantissa x 2^exponent
        fp_value = $itor(result_mantissa) * (2.0 ** $itor(result_exponent));
        
        $display("[TEST] %s", test_name);
        $display("  Inputs: exp_left=%0d, exp_right=%0d", exp_left, exp_right);
        $display("  Output: mantissa=%0d, exponent=%0d", result_mantissa, result_exponent);
        $display("  FP Value: %e (mantissa x 2^%0d)", fp_value, result_exponent);
        $display("");
    endtask
    
    // ===================================================================
    // Test Stimulus
    // ===================================================================
    initial begin
        $display("======================================================");
        $display("  GFP8 Group Dot Product Module Testbench (Registered)");
        $display("======================================================");
        $display("");
        
        // Initialize signals
        reset_n = 0;
        exp_left = 0;
        exp_right = 0;
        man_left = 0;
        man_right = 0;
        
        // Reset sequence
        #20;
        reset_n = 1;
        #20;
        
        // ===============================================================
        // Test 1: Simple known values
        // ===============================================================
        $display("[TEST 1] Simple known values (all 1s)");
        exp_left = 5'd15;   // Bias value
        exp_right = 5'd15;  // Bias value
        
        // All mantissas = 1
        for (int i = 0; i < 32; i++) begin
            man_left[i*8 +: 8] = 8'sd1;
            man_right[i*8 +: 8] = 8'sd1;
        end
        
        // Wait for computation + 1 cycle latency
        @(posedge clk);  // Computation happens
        @(posedge clk);  // Result registered
        display_result("All 1s: 32 x (1 x 1) = 32");
        
        // Expected: mantissa = 32, exponent = 15+15-30 = 0
        assert (result_mantissa == 32) else $error("Mantissa mismatch: expected 32, got %0d", result_mantissa);
        assert (result_exponent == 0) else $error("Exponent mismatch: expected 0, got %0d", result_exponent);
        
        // ===============================================================
        // Test 2: Zero exponent (should return zero)
        // ===============================================================
        $display("[TEST 2] Zero exponent");
        exp_left = 5'd0;
        exp_right = 5'd15;
        
        // Mantissas with non-zero values
        for (int i = 0; i < 32; i++) begin
            man_left[i*8 +: 8] = 8'sd10;
            man_right[i*8 +: 8] = 8'sd20;
        end
        
        // Wait for computation + 1 cycle latency
        @(posedge clk);
        @(posedge clk);
        display_result("Zero exponent -> zero result");
        
        // Expected: mantissa = 0, exponent = 0
        assert (result_mantissa == 0) else $error("Mantissa should be 0, got %0d", result_mantissa);
        assert (result_exponent == 0) else $error("Exponent should be 0, got %0d", result_exponent);
        
        // ===============================================================
        // Test 3: Negative mantissas
        // ===============================================================
        $display("[TEST 3] Negative mantissas");
        exp_left = 5'd16;
        exp_right = 5'd14;
        
        // Mixed positive and negative
        for (int i = 0; i < 16; i++) begin
            man_left[i*8 +: 8] = 8'sd2;
            man_right[i*8 +: 8] = 8'sd3;
        end
        for (int i = 16; i < 32; i++) begin
            man_left[i*8 +: 8] = -8'sd2;
            man_right[i*8 +: 8] = 8'sd3;
        end
        
        // Wait for computation + 1 cycle latency
        @(posedge clk);
        @(posedge clk);
        display_result("Mixed signs: 16x(2x3) + 16x(-2x3) = 96 - 96 = 0");
        
        // Expected: mantissa = 0 (cancellation), exponent varies
        assert (result_mantissa == 0) else $error("Mantissa should be 0, got %0d", result_mantissa);
        
        // ===============================================================
        // Test 4: Actual hex file data (first line)
        // ===============================================================
        $display("[TEST 4] Actual data from left.hex/right.hex (NV 0, Group 0)");
        
        exp_left = 5'd6;   // First exponent from left.hex
        exp_right = 5'd7;  // First exponent from right.hex
        
        // Example mantissa values (pack directly into 256-bit vectors)
        // First 8 elements
        man_left[7:0]     = 8'sd99;  man_right[7:0]     = 8'sd86;
        man_left[15:8]    = 8'sd52;  man_right[15:8]    = 8'sd70;
        man_left[23:16]   = -8'sd74; man_right[23:16]   = 8'sd39;
        man_left[31:24]   = -8'sd58; man_right[31:24]   = -8'sd49;
        man_left[39:32]   = -8'sd7;  man_right[39:32]   = 8'sd19;
        man_left[47:40]   = 8'sd84;  man_right[47:40]   = 8'sd3;
        man_left[55:48]   = 8'sd34;  man_right[55:48]   = 8'sd25;
        man_left[63:56]   = 8'sd29;  man_right[63:56]   = 8'sd30;
        
        // Next 8 elements
        man_left[71:64]   = 8'sd37;  man_right[71:64]   = 8'sd28;
        man_left[79:72]   = 8'sd7;   man_right[79:72]   = -8'sd35;
        man_left[87:80]   = -8'sd40; man_right[87:80]   = -8'sd15;
        man_left[95:88]   = 8'sd51;  man_right[95:88]   = -8'sd51;
        man_left[103:96]  = 8'sd50;  man_right[103:96]  = -8'sd44;
        man_left[111:104] = -8'sd10; man_right[111:104] = 8'sd23;
        man_left[119:112] = 8'sd74;  man_right[119:112] = -8'sd28;
        man_left[127:120] = 8'sd23;  man_right[127:120] = -8'sd18;
        
        // Next 8 elements
        man_left[135:128] = -8'sd41; man_right[135:128] = 8'sd21;
        man_left[143:136] = 8'sd8;   man_right[143:136] = -8'sd12;
        man_left[151:144] = 8'sd24;  man_right[151:144] = 8'sd17;
        man_left[159:152] = -8'sd5;  man_right[159:152] = 8'sd10;
        man_left[167:160] = -8'sd61; man_right[167:160] = 8'sd22;
        man_left[175:168] = -8'sd12; man_right[175:168] = 8'sd28;
        man_left[183:176] = 8'sd61;  man_right[183:176] = 8'sd24;
        man_left[191:184] = -8'sd30; man_right[191:184] = -8'sd15;
        
        // Last 8 elements
        man_left[199:192] = 8'sd2;   man_right[199:192] = 8'sd31;
        man_left[207:200] = -8'sd72; man_right[207:200] = -8'sd23;
        man_left[215:208] = 8'sd23;  man_right[215:208] = 8'sd32;
        man_left[223:216] = -8'sd24; man_right[223:216] = 8'sd30;
        man_left[231:224] = 8'sd78;  man_right[231:224] = -8'sd40;
        man_left[239:232] = -8'sd28; man_right[239:232] = -8'sd34;
        man_left[247:240] = 8'sd47;  man_right[247:240] = -8'sd18;
        man_left[255:248] = 8'sd39;  man_right[255:248] = 8'sd40;
        
        // Wait for computation + 1 cycle latency
        @(posedge clk);
        @(posedge clk);
        display_result("Real data from hex files");
        
        $display("  Manual verification:");
        $display("  - Expected mantissa: sum of 32 products");
        $display("  - Expected exponent: 6 + 7 - 30 = -17");
        
        // ===============================================================
        // Test Complete
        // ===============================================================
        $display("======================================================");
        $display("  All tests completed!");
        $display("======================================================");
        
        #20;
        $finish;
    end

endmodule
