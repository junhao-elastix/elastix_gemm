// ------------------------------------------------------------------
// GFP8 BCV Loop Controller
//
// Purpose: Orchestrate BxCxV nested loops for matrix multiplication
// Algorithm: For each (b,c): accumulate V Native Vector dot products
//
// Matrix Dimensions:
//  - Matrix A (left): B rows x (128xV) columns -> uses BxV Native Vectors
//  - Matrix B (right): (128xV) rows x C columns -> uses CxV Native Vectors
//  - Output: B x C results (one per (b,c) pair)
//
// State Machine:
//  IDLE         -> Wait for TILE command
//  FILL_BUFFER  -> Load complete NV for both NV_left and NV_right (1 cycle)
//                  Direct combinational read from tile_bram's NV interface
//  COMPUTE_NV   -> Compute NV dot product (4 cycles)  
//  ACCUM        -> Accumulate result into V-loop accumulator (1 cycle)
//  RETURN       -> Output final result after V iterations complete (1 cycle)
//
// Latency per output: 6 (pipelined fill) + 4 (compute) + 1 (accum) = 11 cycles per V
//                     Total: 11xV + 1 (return) cycles per BxC result
//                     (Extra 5 cycles per V for 200-300 MHz timing optimization)
//
// OPTIMIZATION: Single-cycle NV read via tile_bram's NV interface
//
// Author: Refactoring from compute_engine.sv
// Date: Fri Oct 10 2025
// ------------------------------------------------------------------

module gfp8_bcv_controller (
    // Clock and Reset
    input  logic        i_clk,
    input  logic        i_reset_n,
    
    // TILE Command Interface
    input  logic        i_tile_en,
    input  logic [7:0]  i_dim_b,              // Output rows (batch)
    input  logic [7:0]  i_dim_c,              // Output columns
    input  logic [7:0]  i_dim_v,              // Inner dimension multiplier (V Native Vectors)
    input  logic [8:0]  i_left_base_addr,     // Base address for left matrix in tile_bram (9-bit for 512 lines)
    input  logic [8:0]  i_right_base_addr,    // Base address for right matrix in tile_bram (9-bit for 512 lines)
    output logic        o_tile_done,

    // Native Vector Read Interface (to tile_bram)
    output logic [6:0]   o_nv_left_rd_idx,      // NV index [0-127]
    input  logic [31:0]  i_nv_left_exp,         // Packed exponents
    input  logic [255:0] i_nv_left_man [0:3],   // 4 mantissa groups
    
    output logic [6:0]   o_nv_right_rd_idx,     // NV index [0-127]
    input  logic [31:0]  i_nv_right_exp,        // Packed exponents
    input  logic [255:0] i_nv_right_man [0:3],  // 4 mantissa groups
    
    // Result Interface
    output logic signed [31:0] o_result_mantissa,
    output logic signed [7:0]  o_result_exponent,
    output logic               o_result_valid
);

    // ===================================================================
    // State Machine Definition
    // ===================================================================
    typedef enum logic [2:0] {
        ST_IDLE        = 3'd0,
        ST_FILL_BUFFER = 3'd1,  // Load both NV_left and NV_right (4 cycles)
        ST_COMPUTE_NV  = 3'd2,  // Compute NV dot product (2 cycles)
        ST_ACCUM       = 3'd3,  // Accumulate into V-loop accumulator
        ST_RETURN      = 3'd4,  // Output final result
        ST_DONE        = 3'd5
    } state_t;
    
    state_t state_reg, state_next;
    
    // ===================================================================
    // Loop Indices (B, C, V nested loops)
    // ===================================================================
    logic [7:0] b_idx;  // Batch index (0 to B-1)
    logic [7:0] c_idx;  // Column index (0 to C-1)
    logic [7:0] v_idx;  // Vector index (0 to V-1)
    
    // Dimension registers
    logic [7:0] dim_b_reg, dim_c_reg, dim_v_reg;
    logic [8:0] left_base_reg, right_base_reg;  // 9-bit for 512-line tile_bram
    
    // Rising edge detection for i_tile_en
    logic i_tile_en_prev;
    logic i_tile_en_rising;
    
    assign i_tile_en_rising = i_tile_en && !i_tile_en_prev;
    
    // Fill buffer ready flag (set when last group captured)
    logic fill_buffer_ready;
    
    // ===================================================================
    // Native Vector Buffers (Local Storage)
    // ===================================================================
    
    // NV_left buffer
    logic [31:0]  nv_left_exp;         // 4 bytes (one per group)
    logic [255:0] nv_left_man [0:3];   // 4 lines x 256 bits
    
    // NV_right buffer
    logic [31:0]  nv_right_exp;        // 4 bytes (one per group)
    logic [255:0] nv_right_man [0:3];  // 4 lines x 256 bits
    
    // No fill cycle counter needed - single-cycle NV read
    
    // ===================================================================
    // NV Dot Product Instance
    // ===================================================================
    logic signed [31:0] nv_dot_mantissa;
    logic signed [7:0]  nv_dot_exponent;
    
    // Enable signal: pulse high when entering ST_COMPUTE_NV
    logic nv_dot_input_valid;
    assign nv_dot_input_valid = (state_reg != ST_COMPUTE_NV) && (state_next == ST_COMPUTE_NV);
    
    gfp8_nv_dot u_nv_dot (
        .i_clk              (i_clk),
        .i_reset_n          (i_reset_n),
        .i_input_valid      (nv_dot_input_valid),  // Latch inputs only when entering COMPUTE
        .i_exp_left         (nv_left_exp),
        .i_man_left         (nv_left_man),
        .i_exp_right        (nv_right_exp),
        .i_man_right        (nv_right_man),
        .o_result_mantissa  (nv_dot_mantissa),
        .o_result_exponent  (nv_dot_exponent)
    );
    
    // ===================================================================
    // V-Loop Accumulator
    // ===================================================================
    logic signed [31:0] accum_mantissa;
    logic signed [7:0]  accum_exponent;
    
    // Compute pipeline counter (track 4-cycle latency)
    logic [2:0] compute_wait;
    
    // ===================================================================
    // State Machine - Next State Logic
    // ===================================================================
    always_comb begin
        state_next = state_reg;
        
        case (state_reg)
            ST_IDLE: begin
                if (i_tile_en_rising) begin
                    state_next = ST_FILL_BUFFER;
                end
            end
            
            ST_FILL_BUFFER: begin
                // Wait for NV data to be latched before transitioning
                if (fill_buffer_ready) begin
                    state_next = ST_COMPUTE_NV;
                end
            end
            
            ST_COMPUTE_NV: begin
                // Wait for gfp8_nv_dot 4-cycle pipeline
                if (compute_wait == 3'd3) begin
                    state_next = ST_ACCUM;
                end
            end
            
            ST_ACCUM: begin
                // Check if V loop is complete
                if (v_idx >= dim_v_reg - 1) begin
                    state_next = ST_RETURN;
                end else begin
                    // More V iterations needed
                    state_next = ST_FILL_BUFFER;
                end
            end
            
            ST_RETURN: begin
                // Check if all BxC outputs are complete
                if (c_idx >= dim_c_reg - 1 && b_idx >= dim_b_reg - 1) begin
                    state_next = ST_DONE;
                end else begin
                    // Start next output element (next b,c pair)
                    state_next = ST_FILL_BUFFER;
                end
            end
            
            ST_DONE: begin
                state_next = ST_IDLE;
            end
            
            default: state_next = ST_IDLE;
        endcase
    end
    
    // ===================================================================
    // State Machine - Sequential Logic
    // ===================================================================
    always_ff @(posedge i_clk or negedge i_reset_n) begin
        if (!i_reset_n) begin
            state_reg <= ST_IDLE;
        end else begin
            state_reg <= state_next;
        end
    end
    
    // ===================================================================
    // NV Read Index Generation - PIPELINED for 200-300 MHz (TIMING OPTIMIZATION)
    // ===================================================================
    // Add pipeline register to break critical path:
    // Before: v_idx → index_calc → tile_bram (8.5ns - too long!)
    // After:  v_idx → index_calc → INDEX_REG → tile_bram (split into 2 stages)
    
    // Combinational NV index calculation
    logic [6:0] left_nv_index_comb, right_nv_index_comb;
    logic [6:0] left_base_nv, right_base_nv;
    
    // Convert base addresses from line units to NV units (divide by 4)
    assign left_base_nv = left_base_reg[8:2];
    assign right_base_nv = right_base_reg[8:2];
    
    always_comb begin
        // Calculate NV indices combinationally
        left_nv_index_comb = left_base_nv + (b_idx * dim_v_reg + v_idx);
        right_nv_index_comb = right_base_nv + (c_idx * dim_v_reg + v_idx);
    end
    
    // PIPELINE REGISTER: Break timing path here
    logic [6:0] left_nv_index_reg, right_nv_index_reg;
    logic       nv_indices_valid;
    
    always_ff @(posedge i_clk or negedge i_reset_n) begin
        if (!i_reset_n) begin
            left_nv_index_reg <= 7'd0;
            right_nv_index_reg <= 7'd0;
            nv_indices_valid <= 1'b0;
        end else begin
            // Register indices during FILL_BUFFER state
            if (state_reg == ST_FILL_BUFFER && !fill_buffer_ready) begin
                left_nv_index_reg <= left_nv_index_comb;
                right_nv_index_reg <= right_nv_index_comb;
                nv_indices_valid <= 1'b1;
                `ifdef SIMULATION
                $display("[NV_IDX] @%0t Registered Left NV[%0d], Right NV[%0d] for B=%0d, C=%0d, V=%0d", 
                         $time, left_nv_index_comb, right_nv_index_comb, b_idx, c_idx, v_idx);
                `endif
            end else if (state_reg != ST_FILL_BUFFER) begin
                nv_indices_valid <= 1'b0;
            end
        end
    end
    
    // Output registered indices to tile_bram
    assign o_nv_left_rd_idx = left_nv_index_reg;
    assign o_nv_right_rd_idx = right_nv_index_reg;
    
    // ===================================================================
    // Buffer Filling Logic (Single-cycle NV capture)
    // ===================================================================
    always_ff @(posedge i_clk or negedge i_reset_n) begin
        if (!i_reset_n) begin
            fill_buffer_ready <= 1'b0;
            nv_left_exp <= 32'd0;
            nv_right_exp <= 32'd0;
            for (int i = 0; i < 4; i++) begin
                nv_left_man[i] <= 256'd0;
                nv_right_man[i] <= 256'd0;
            end
        end else begin
            case (state_reg)
                ST_IDLE: begin
                    fill_buffer_ready <= 1'b0;
                end
                
                ST_FILL_BUFFER: begin
                    // PIPELINED: Cycle 0 = calc indices, Cycle 1 = wait for BRAM, Cycles 2-5 = capture groups
                    if (fill_cycle == 3'd1 && nv_indices_valid) begin
                        // Cycle 1: Indices now registered, start BRAM read for G0
                        // BRAM data will be ready next cycle
                    end else if (fill_cycle == 3'd2) begin
                        // Cycle 2: Capture G0 (from previous cycle's read)
                        nv_left_exp[7:0] <= i_nv_left_exp[7:0];
                        nv_right_exp[7:0] <= i_nv_right_exp[7:0];
                        nv_left_man[0] <= i_nv_left_man[0];
                        nv_right_man[0] <= i_nv_right_man[0];
                    end else if (fill_cycle == 3'd3) begin
                        // Cycle 3: Capture G1
                        nv_left_exp[15:8] <= i_nv_left_exp[15:8];
                        nv_right_exp[15:8] <= i_nv_right_exp[15:8];
                        nv_left_man[1] <= i_nv_left_man[1];
                        nv_right_man[1] <= i_nv_right_man[1];
                    end else if (fill_cycle == 3'd4) begin
                        // Cycle 4: Capture G2
                        nv_left_exp[23:16] <= i_nv_left_exp[23:16];
                        nv_right_exp[23:16] <= i_nv_right_exp[23:16];
                        nv_left_man[2] <= i_nv_left_man[2];
                        nv_right_man[2] <= i_nv_right_man[2];
                    end else if (fill_cycle == 3'd5) begin
                        // Cycle 5: Capture G3 and set ready flag
                        nv_left_exp[31:24] <= i_nv_left_exp[31:24];
                        nv_right_exp[31:24] <= i_nv_right_exp[31:24];
                        nv_left_man[3] <= i_nv_left_man[3];
                        nv_right_man[3] <= i_nv_right_man[3];
                        fill_buffer_ready <= 1'b1;
                        `ifdef SIMULATION
                        $display("[BCV_FILL] @%0t Captured all 4 groups for B=%0d, C=%0d, V=%0d (PIPELINED)",
                                 $time, b_idx, c_idx, v_idx);
                        $display("  Left exp: 0x%08x, Right exp: 0x%08x", {i_nv_left_exp[31:24], nv_left_exp[23:0]}, {i_nv_right_exp[31:24], nv_right_exp[23:0]});
                        `endif
                    end
                    
                    // Increment fill cycle counter
                    if (fill_cycle < 3'd5) begin
                        fill_cycle <= fill_cycle + 1;
                    end else if (fill_buffer_ready) begin
                        fill_cycle <= 3'd0;  // Reset after ready
                    end
                end
                
                ST_COMPUTE_NV: begin
                    // Clear the ready flag once we've transitioned
                    fill_buffer_ready <= 1'b0;
                end
                
                default: begin
                    // Keep default values
                end
            endcase
        end
    end
    
    // ===================================================================
    // Compute Pipeline Control
    // ===================================================================
    always_ff @(posedge i_clk or negedge i_reset_n) begin
        if (!i_reset_n) begin
            compute_wait <= 3'd0;
        end else begin
            case (state_reg)
                ST_COMPUTE_NV: begin
                    if (compute_wait < 3'd3) begin
                        compute_wait <= compute_wait + 1;  // Count: 0→1→2→3
                    end
                end
                default: begin
                    compute_wait <= 3'd0;
                end
            endcase
        end
    end
    
    // ===================================================================
    // V-Loop Accumulation (with Exponent Alignment)
    // ===================================================================
    always_ff @(posedge i_clk or negedge i_reset_n) begin
        if (!i_reset_n) begin
            accum_mantissa <= 32'sd0;
            accum_exponent <= 8'sd0;
        end else begin
            case (state_reg)
                ST_IDLE: begin
                    accum_mantissa <= 32'sd0;
                    accum_exponent <= 8'sd0;
                end
                
                ST_ACCUM: begin
                    if (v_idx == 8'd0) begin
                        // First V iteration - initialize accumulator
                        accum_mantissa <= nv_dot_mantissa;
                        accum_exponent <= nv_dot_exponent;
                        `ifdef SIMULATION
                        $display("[BCV_ACCUM] @%0t [B%0d,C%0d] V=%0d INIT: mant=%0d (0x%08x), exp=%0d",
                                 $time, b_idx, c_idx, v_idx, nv_dot_mantissa, nv_dot_mantissa, nv_dot_exponent);
                        `endif
                    end else begin
                        // Accumulate with exponent alignment (FIXED: match original implementation)
                        automatic logic signed [7:0] max_exp;
                        automatic logic [7:0] exp_diff_accum, exp_diff_dot;
                        automatic logic signed [31:0] aligned_accum, aligned_dot;
                        automatic logic signed [31:0] sum_mantissa;
                        
                        // Find maximum exponent (using signed comparison for negative exponents)
                        if ($signed(accum_exponent) > $signed(nv_dot_exponent)) begin
                            max_exp = accum_exponent;
                        end else begin
                            max_exp = nv_dot_exponent;
                        end
                        
                        // Align mantissas to maximum exponent
                        exp_diff_accum = max_exp - accum_exponent;
                        exp_diff_dot = max_exp - nv_dot_exponent;
                        
                        // Align accumulated mantissa with underflow check
                        if (exp_diff_accum > 31) begin
                            aligned_accum = 32'sd0;  // Underflow - set to zero
                        end else begin
                            aligned_accum = $signed(accum_mantissa) >>> exp_diff_accum;
                        end
                        
                        // Align dot product mantissa with underflow check
                        if (exp_diff_dot > 31) begin
                            aligned_dot = 32'sd0;  // Underflow - set to zero
                        end else begin
                            aligned_dot = $signed(nv_dot_mantissa) >>> exp_diff_dot;
                        end
                        
                        // Sum aligned mantissas
                        sum_mantissa = aligned_accum + aligned_dot;
                        
                        // Update accumulator
                        accum_mantissa <= sum_mantissa;
                        accum_exponent <= max_exp;
                        `ifdef SIMULATION
                        $display("[BCV_ACCUM] @%0t [B%0d,C%0d] V=%0d ADD: accum_m=%0d(exp=%0d), dot_m=%0d(exp=%0d) -> aligned_a=%0d, aligned_d=%0d -> sum=%0d(exp=%0d)",
                                 $time, b_idx, c_idx, v_idx, accum_mantissa, accum_exponent, nv_dot_mantissa, nv_dot_exponent,
                                 aligned_accum, aligned_dot, sum_mantissa, max_exp);
                        `endif
                    end
                end
                
                ST_RETURN: begin
                    // Reset accumulator for next BxC output (after outputting result)
                    accum_mantissa <= 32'sd0;
                    accum_exponent <= 8'sd0;
                end
            endcase
        end
    end
    
    // ===================================================================
    // Loop Index Control (B, C, V nested loops)
    // ===================================================================
    always_ff @(posedge i_clk or negedge i_reset_n) begin
        if (!i_reset_n) begin
            b_idx <= 8'd0;
            c_idx <= 8'd0;
            v_idx <= 8'd0;
            dim_b_reg <= 8'd0;
            dim_c_reg <= 8'd0;
            dim_v_reg <= 8'd0;
            left_base_reg <= 11'd0;
            right_base_reg <= 11'd0;
            i_tile_en_prev <= 1'b0;
        end else begin
            // Update previous value for edge detection
            i_tile_en_prev <= i_tile_en;
            
            case (state_reg)
                ST_IDLE: begin
                    if (i_tile_en_rising) begin
                        // Capture dimensions
                        dim_b_reg <= i_dim_b;
                        dim_c_reg <= i_dim_c;
                        dim_v_reg <= i_dim_v;
                        left_base_reg <= i_left_base_addr;
                        right_base_reg <= i_right_base_addr;
                        // Initialize indices
                        b_idx <= 8'd0;
                        c_idx <= 8'd0;
                        v_idx <= 8'd0;
                        $display("[BCV_LOOP] @%0t NEW TILE: B=%0d, C=%0d, V=%0d, left_base=%0d, right_base=%0d", 
                                 $time, i_dim_b, i_dim_c, i_dim_v, i_left_base_addr, i_right_base_addr);
                        $display("[BCV_LOOP] @%0t DIM_CAPTURE: dim_b_reg=%0d->%0d, dim_c_reg=%0d->%0d, dim_v_reg=%0d->%0d",
                                 $time, dim_b_reg, i_dim_b, dim_c_reg, i_dim_c, dim_v_reg, i_dim_v);
                    end
                end
                
                ST_ACCUM: begin
                    // Check if V loop is complete before advancing
                    if (v_idx < dim_v_reg - 1) begin
                        // More V iterations needed - advance V index
                        v_idx <= v_idx + 1;
                        $display("[BCV_LOOP] ACCUM: b=%0d, c=%0d, v=%0d -> v=%0d", 
                                 b_idx, c_idx, v_idx, v_idx + 1);
                    end
                    // If v_idx >= dim_v_reg - 1, don't increment (going to RETURN state)
                end
                
                ST_RETURN: begin
                    // V loop complete, advance C and B indices
                    v_idx <= 8'd0;  // Reset V for next (b,c) pair
                    
                    $display("[BCV_LOOP] RETURN: b=%0d, c=%0d completed V loop, advancing indices", 
                             b_idx, c_idx);
                    
                    // Only advance indices if NOT done with all outputs
                    if (!(c_idx >= dim_c_reg - 1 && b_idx >= dim_b_reg - 1)) begin
                        // Advance C index
                        if (c_idx >= dim_c_reg - 1) begin
                            c_idx <= 8'd0;
                            // Advance B index
                            b_idx <= b_idx + 1;
                            $display("[BCV_LOOP]   -> Next: b=%0d, c=0", b_idx + 1);
                        end else begin
                            c_idx <= c_idx + 1;
                            $display("[BCV_LOOP]   -> Next: b=%0d, c=%0d", b_idx, c_idx + 1);
                        end
                    end else begin
                        $display("[BCV_LOOP]   -> DONE (all BxC outputs complete)");
                    end
                end
            endcase
        end
    end
    
    // ===================================================================
    // Output Control
    // ===================================================================
    always_ff @(posedge i_clk or negedge i_reset_n) begin
        if (!i_reset_n) begin
            o_result_mantissa <= 32'sd0;
            o_result_exponent <= 8'sd0;
            o_result_valid <= 1'b0;
            o_tile_done <= 1'b0;
        end else begin
            // Default
            o_result_valid <= 1'b0;
            o_tile_done <= 1'b0;
            
            case (state_reg)
                ST_RETURN: begin
                    // Output accumulated result for this (b,c) pair
                    o_result_mantissa <= accum_mantissa;
                    o_result_exponent <= accum_exponent;
                    o_result_valid <= 1'b1;
                    `ifdef SIMULATION
                    $display("[BCV_ACCUM] @%0t [B%0d,C%0d] RETURN: Final GFP result = mant=%0d (0x%08x), exp=%0d",
                             $time, b_idx, c_idx, accum_mantissa, accum_mantissa, accum_exponent);
                    `endif
                end
                
                ST_DONE: begin
                    o_tile_done <= 1'b1;
                end
            endcase
        end
    end

endmodule

